// 1.14 inch 240x135 SPI LCD TEST for TANG NANO 9K
// by fanoble, QQ:87430545
// 27/6/2022

`timescale 1ps/1ps

module lcd114_test(
	input clk, // 27M
	input resetn,

	output ser_tx,
	input ser_rx,

	output lcd_resetn,
	output lcd_clk,
	output lcd_cs,
	output lcd_rs,
	output lcd_data
);

localparam MAX_CMDS = 69;

wire [8:0] init_cmd[MAX_CMDS:0];

assign init_cmd[ 0] = 9'h036;
assign init_cmd[ 1] = 9'h170;
assign init_cmd[ 2] = 9'h03A;
assign init_cmd[ 3] = 9'h105;
assign init_cmd[ 4] = 9'h0B2;
assign init_cmd[ 5] = 9'h10C;
assign init_cmd[ 6] = 9'h10C;
assign init_cmd[ 7] = 9'h100;
assign init_cmd[ 8] = 9'h133;
assign init_cmd[ 9] = 9'h133;
assign init_cmd[10] = 9'h0B7;
assign init_cmd[11] = 9'h135;
assign init_cmd[12] = 9'h0BB;
assign init_cmd[13] = 9'h119;
assign init_cmd[14] = 9'h0C0;
assign init_cmd[15] = 9'h12C;
assign init_cmd[16] = 9'h0C2;
assign init_cmd[17] = 9'h101;
assign init_cmd[18] = 9'h0C3;
assign init_cmd[19] = 9'h112;
assign init_cmd[20] = 9'h0C4;
assign init_cmd[21] = 9'h120;
assign init_cmd[22] = 9'h0C6;
assign init_cmd[23] = 9'h10F;
assign init_cmd[24] = 9'h0D0;
assign init_cmd[25] = 9'h1A4;
assign init_cmd[26] = 9'h1A1;
assign init_cmd[27] = 9'h0E0;
assign init_cmd[28] = 9'h1D0;
assign init_cmd[29] = 9'h104;
assign init_cmd[30] = 9'h10D;
assign init_cmd[31] = 9'h111;
assign init_cmd[32] = 9'h113;
assign init_cmd[33] = 9'h12B;
assign init_cmd[34] = 9'h13F;
assign init_cmd[35] = 9'h154;
assign init_cmd[36] = 9'h14C;
assign init_cmd[37] = 9'h118;
assign init_cmd[38] = 9'h10D;
assign init_cmd[39] = 9'h10B;
assign init_cmd[40] = 9'h11F;
assign init_cmd[41] = 9'h123;
assign init_cmd[42] = 9'h0E1;
assign init_cmd[43] = 9'h1D0;
assign init_cmd[44] = 9'h104;
assign init_cmd[45] = 9'h10C;
assign init_cmd[46] = 9'h111;
assign init_cmd[47] = 9'h113;
assign init_cmd[48] = 9'h12C;
assign init_cmd[49] = 9'h13F;
assign init_cmd[50] = 9'h144;
assign init_cmd[51] = 9'h151;
assign init_cmd[52] = 9'h12F;
assign init_cmd[53] = 9'h11F;
assign init_cmd[54] = 9'h11F;
assign init_cmd[55] = 9'h120;
assign init_cmd[56] = 9'h123;
assign init_cmd[57] = 9'h021;
assign init_cmd[58] = 9'h029;

assign init_cmd[59] = 9'h02A; // column
assign init_cmd[60] = 9'h100;
assign init_cmd[61] = 9'h128;
assign init_cmd[62] = 9'h101;
assign init_cmd[63] = 9'h117;
assign init_cmd[64] = 9'h02B; // row
assign init_cmd[65] = 9'h100;
assign init_cmd[66] = 9'h135;
assign init_cmd[67] = 9'h100;
assign init_cmd[68] = 9'h1BB;
assign init_cmd[69] = 9'h02C; // start

localparam INIT_RESET   = 4'b0000; // delay 100ms while reset
localparam INIT_PREPARE = 4'b0001; // delay 200ms after reset
localparam INIT_WAKEUP  = 4'b0010; // write cmd 0x11 MIPI_DCS_EXIT_SLEEP_MODE
localparam INIT_SNOOZE  = 4'b0011; // delay 120ms after wakeup
localparam INIT_WORKING = 4'b0100; // write command & data
localparam INIT_DONE    = 4'b0101; // all done

`ifdef MODELTECH

localparam CNT_100MS = 32'd2700000;
localparam CNT_120MS = 32'd3240000;
localparam CNT_200MS = 32'd5400000;

`else

// speedup for simulation
localparam CNT_100MS = 32'd27;
localparam CNT_120MS = 32'd32;
localparam CNT_200MS = 32'd54;

`endif


reg [ 3:0] init_state;
reg [ 6:0] cmd_index;
reg [31:0] clk_cnt;
reg [ 4:0] bit_loop;

reg [15:0] pixel_cnt;

reg lcd_cs_r;
reg lcd_rs_r;
reg lcd_reset_r;

reg [7:0] spi_data;

assign lcd_resetn = lcd_reset_r;
assign lcd_clk    = ~clk;
assign lcd_cs     = lcd_cs_r;
assign lcd_rs     = lcd_rs_r;
assign lcd_data   = spi_data[7]; // MSB

// gen color bar
//wire [15:0] pixel = (pixel_cnt >= 21600) ? 16'h0000 :
//					(pixel_cnt >= 10800) ? 16'hffff : 16'heeee;
reg [3:0] time_cnt;
wire [32399:0]cxk[9:0];
assign cxk[0][32399:0] = 32400'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003e0000000000000000000000000000000000000000000000000000000003ffc00000000000000000000000000000000000000000000000000000000ffff00000000000000000000000000000000000000000000000000000001fffff0000000000000000000000000000000000000000000000000000007fffffffc000000000000000000000000000000000000000000000000001ffffffffe000000000000000000000000000000000000000000000000007fffffffff800000000000000000000000000000000000000000000000007fffffffffc0000000000000000000000000000000000000000000000000ffffffffffe0000000000000000000000000000000000000000000000000fffffffffff0000000000000000000000000000000000000000000000001fffffffffff8000000000000000000000000000000000000000000000003fffffffffffc000000000000000000000000000000000000000000000003fffffffffffe000000000000000000000000000000000000000000000003fffffffffffe000000000000000000000000000000000000000000000003fffffffffffe000000000000000000000000000000000000000000000003fffffffffffe000000000000000000000000000000000000000000000003fffffffffffe000000000000000000000000000000000000000000000003ffffffffffff000000000000000000000000000000000000000000000003ffffffffffff000000000000000000000000000000000000000000000001ffffffffffff000000000000000000000000000000000000000000000001fffffffffffe000000000000000000000000000000000000000000000001fffffffffffe000000000000000000000000000000000000000000000001fffffffffffe000000000000000000000000000000000000000000000000fffffffffffc000000000000000000000000000000000000000000000000fffffffffff8000000000000000000000000000000000000000000000000fffffffffff8000000000000000000000000000000000000000000000000fffffffffff0000000000000000000000000000000000000000000000000ffffffffffe0000000000000000000000000000000000000000000000000ffffffffff80000000000000000000000000000000000000000000000003ffffffffff8000000000000000000000000000000000000000000000003fffffffffff000000000000000000000000000000000000000000000001ffffffffffff000000000000000000000000000000000000000000000007fffffffffffe00000000000000000000000000000000000000000000001ffffffffffffc0000000000000000000000000000000000000000000007fffffffffffffc000000000000000000000000000000000000000000003ffffffffffffffc00000000000000000000000000000000000000000000fffffffffffffffc00000000000000000000000000000000000000000007fffffffffffffffe0000000000000000000000000000000000000000003ffffffffffffffffe000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000000000000000000007ffffffffffffffffff00000000000000000000000000000000000000007fffffffffffffffffff8000000000000000000000000000000000000001ffffffffffffffffffffc000000000000000000000000000000000000007ffffffffffffffffffffe00000000000000000000000000000000000001ffffffffffffffffffffff00000000000000000000000000000000000007ffffffffffffffffffffff8000000000000000000000000000000000000fffffffffffffffffffffffc000000000000000000000000000000000001fffffffffffffffffffffffc000000000000000000000000000000000007fffffffffffffffffffffffe00000000000000000000000000000000000fffffffffffffffffffffffff00000000000000000000000000000000001fffffffffffffffffffffffff80000000000000000000000000000000003fffffffffffffffffffffffffc000000000000000000000000000000000ffffffffffffffffffffffffffe000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000007ffffffffffffffffffffffffffc00000000000000000000000000000001fffffffffffffffffffffffffffc00000000000000000000000000000003fffffffffffffffffffffffffffc00000000000000000000000000000007fffffffffffffffffffffffffffc0000000000000000000000000000001ffffffffffffffffffffffffffffc0000000000000000000000000000007ffffffffffffffffffffffffffff8000000000000000000000000000000fffffffffffffffffffffffffffff8000000000000000000000000000003fffffffffffffffffffffffffffff8000000000000000000000000000007fffffffffffffffffffffffffffff8000000000000000000000000000007fffffffffffffffffffffffffffff800000000000000000000000000000ffffffffffffffffffffffffffffff800000000000000000000000000000fffff80fffffffffffffffffffffff800000000000000000000000000001ffffc007ffffffffffffffffffffff000000000000000000000000000001ffffc003ffffffffffffffffffffff000000000000000000000000000001ffff8003ffffffffffffffffffffff000000000000000000000000000001ffff8003ffffffffffffffffffffff000000000000000000000000000001ffff8003ffffffffffffffffffffff000000000000000000000000000000ffff8003ffffffffffffffffffffff000000000000000000000000000000ffff8007ffffffffffffffffffffff0000000000000000000000000000007fffc007fffffffffffffffffffffe0000000000000000000000000000007fffc00ffffffffffffffffffffffe0000000000000000000000000000003fffe01ffffffffffffffffffffffe0000000000000000000000000000001ffffffffffffffffffffffffffffe0000000000000000000000000000001ffffffffffffffffffffffffffffc0000000000000000000000000000000ffffffffffffffffffffffffffff800000000000000000000000000000007fffffffffffffffffffffffffff800000000000000000000000000000003fffffffffffffffffffffffffff000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000ff00000000000001ffffffffffffffffffffffffffffc000000000000000ff00000000000001ffffffffffffffffffffffffffff8000000000000000ff00000000000001ffffffffffffffffffffffffffff0000000000000000ff00000000000001ffbfffffffffffffffffffffffff0000000000000000ff000001ff000001ff9ffffffffffffffffffffffffe0000000000000000ff000003ff980001ff8ffffffffffffffffffffffffc0000000000000000ff000007fff80001ff87fffffffffffffffffffffffc0000000000000000ff000007fff80001ff83fffffffffffffffffffffff80000000000000000ff000007fffc0001ff81fffffffffffffffffffffff80000000000000000ff00001ffff00001ff80fffffffffffffffffffffff00000000000000000ff00000fffe00001ff807ffffffffffffffffffffff00000000000000000ff000007ffe00001ff803fffffffffffffffffffffe00000000000000000ff000007ff800001ff803fffffffffffffffffffffc00000000000000000ff000007ff800001ff803fffffffffffffffffffffc00000000000000000ff000001ff000001ff803fffffffffffffffffffff800000000000000000ff080000f8000001ff807ffffffffffffffffffffe000000000000000000ff3e0007fe000001ff80fffffffffffffffffffffc000000000000000000ffff800fff800e01ff81fffffffffffffffffffff8000000000000000000ffffc01fffc07f01ff87fffffffffffffffffffff0000000000000000000ffffff3fffe1ff81ff8fffffffffffffffffffffe0000000000000000000ffffffffffffffc1ff9fffffffffffffffffffffc0000000000000000000ffd3ff8fffffffe1ffbfffffffffffffffffffff80000000000000000000ff811c0fffdffff9ffbfffffffffffffffffffff00000000000000000000ff00000fffc040fdfffffffffffffffffffffffe00000000000000000000ff00000fffc0007ffffffffffffffffffffffffc00000000000000000000ff00000ffee00001fffffffffffffffffffffff000000000000000000000ff000007fe400001ffffffffffffffffffffffe000000000000000000000ff000007fe000001ffffffffffffffffffffffe000000000000000000000ff00000fff000001ffffffffffffffffffffffe000000000000000000000ff000007ff000001ffffffffffffffffffffffe000000000000000000000ff00000fff000001ffffffffffffffffffffffe000000000000000000000;
assign cxk[1][32399:0] = 32400'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003c0000000000000000000000000000000000000000000000000000000001ff8000000000000000000000000000000000000000000000000000000007fff00000000000000000000000000000000000000000000000000000001fffff8000000000000000000000000000000000000000000000000000007ffffffc0000000000000000000000000000000000000000000000000000fffffffe0000000000000000000000000000000000000000000000000001ffffffff0000000000000000000000000000000000000000000000000003ffffffff8000000000000000000000000000000000000000000000000007ffffffffe00000000000000000000000000000000000000000000000000ffffffffff00000000000000000000000000000000000000000000000003ffffffffff00000000000000000000000000000000000000000000000003ffffffffff80000000000000000000000000000000000000000000000003ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe0000000000000000000000000000000000000000000000007ffffffffffe000000000000000000000000000000000000000000000000fffffffffffe000000000000000000000000000000000000000000000007fffffffffffe00000000000000000000000000000000000000000000003ffffffffffffc000000000000000000000000000000000000000000003ffffffffffffff800000000000000000000000000000000000000000001fffffffffffffff00000000000000000000000000000000000000000001fffffffffffffffe00000000000000000000000000000000000000000007fffffffffffffffc0000000000000000000000000000000000000000001ffffffffffffffff8000000000000000000000000000000000000000000fffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff00000000000000000000000000000000000000001ffffffffffffffffffe00000000000000000000000000000000000000007ffffffffffffffffffc0000000000000000000000000000000000000000fffffffffffffffffffc0000000000000000000000000000000000000003fffffffffffffffffffc0000000000000000000000000000000000000007fffffffffffffffffffc000000000000000000000000000000000000000ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffe000000000000000000000000000000000000007fffffffffffffffffffff000000000000000000000000000000000000007fffffffffffffffffffff80000000000000000000000000000000000000ffffffffffffffffffffff80000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000007ffffffffffffffffffffffe000000000000000000000000000000000000ffffffffffffffffffffffff000000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffe0000000000000000000000000000000001ffffffffffffffffffffffffff0000000000000000000000000000000007ffffffffffffffffffffffffff000000000000000000000000000000000fffffffffffffffffffffffffff800000000000000000000000000000001fffffffffffffffffffffffffffc00000000000000000000000000000003fffffffffffffffffffffffffffc00000000000000000000000000000007fffffffffffffffffffffffffffe0000000000000000000000000000001ffffff0fffffffffffffffffffffe0000000000000000000000000000003fffffc07ffffffffffffffffffffc0000000000000000000000000000007fffff803ffffffffffffffffffffc000000000000000000000000000000ffffff803ffffffffffffffffffffc000000000000000000000000000001ffffff003ffffffffffffffffffffc000000000000000000000000000007fffffe003ffffffffffffffffffffc00000000000000000000000000000ffffffc003ffffffffffffffffffffc00000000000000000000000000000ffffff8003ffffffffffffffffffffc00000000000000000000000000001ffffff0003ffffffffffffffffffffc00000000000000000000000000001fffffe0003ffffffffffffffffffffc00000000000000000000000000003fffffe0003ffffffffffffffffffffc00000000000000000000000000003fffffc0003ffffffffffffffffffffc00000000000000000000000000001fffffc0007ffffffffffffffffffffe00000000000000000000000000000fffffc0007ffffffffffffffffffffe000000000000000000000000000007ffffc0007ffffffffffffffffffffe000000000000000000000000000003ffffc000ffffffffffffffffffffff000000000000000000000000000003ffffc001ffffffffffffffffffffff000000000000000000000000000000ffffe001ffffffffffffffffffffff0000000000000000000000000000007ffff003ffffffffffffffffffffff8000000000000000000000000000003ffff807ffffffffffffffffffffff8000000000000000000000000000000ffffc0fffffffffffffffffffffff80000000000000000000000000000007ffffffffffffffffffffffffffff80000000000000000000000000000003ffffffffffffffffffffffffffff80000000000000000000000000000001ffffffffffffffffffffffffffff800000000000000000000000000000007fffffffffffffffffffffffffff800000000000000000000000000000003fffffffffffffffffffffffffff800000000000000000000000000000001fffffffffffffffffffffffffff000000000000000000000000000000000fffffffffffffffffffffffffff0000000000000000000000000000000003fffffffffffffffffffffffffe0000000000000000000000000000000001fffffffffffffffffffffffffe00000000000000000000000000000000007ffffffffffffffffffffffffe00000000000000000000000000000000003ffffffffffffffffffffffffe00000000000000000000000000000000000ffffffffffffffffffffffffc000000000000000000000000000000000007fffffffffffffffffffffff8000000000000000000000000000000000003fffffffffffffffffffffff0000000000000000000000000000000000000fffffffffffffffffffffff00000000000000000000000000000000000007ffffffffffffffffffffff000000000000000000ff00000000000001ff87fffffffffffffffffffffe000000000000000000ff00000000000001ff83fffffffffffffffffffffe000000000000000000ff00000000000001ff83fffffffffffffffffffffe000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff000001ff000001ff83fffffffffffffffffffffc000000000000000000ff000003ff980001ff83fffffffffffffffffffffc000000000000000000ff000007fff80001ff83fffffffffffffffffffff8000000000000000000ff000007fff80001ff8ffffffffffffffffffffff0000000000000000000ff000007fffc0001ff9ffffffffffffffffffffff0000000000000000000ff00001ffff00001ffffffffffffffffffffffffc0000000000000000000ff00000fffe00001ffffffffffffffffffffffff80000000000000000000ff000007ffe00001fffffffffffffffffffffffe00000000000000000000ff000007ff800001ffffffffffffffffffffff0000000000000000000000ff000007ff800001fffffffffffffffffffffc0000000000000000000000ff000001ff000001fffffffffffffffffffff80000000000000000000000ff080000f8000001fffffffffffffffffffff80000000000000000000000ff3e0007fe000001fffffffffffffffffffff80000000000000000000000ffff800fff800e01fffffffffffffffffffff80000000000000000000000ffffc01fffc07f01fffffffffffffffffffff80000000000000000000000ffffff3fffe1ff81fffffffffffffffffffffc0000000000000000000000ffffffffffffffc1fffffffffffffffffffffc0000000000000000000000ff93ff8fffffffe1fffffffffffffffffffffc0000000000000000000000ff811c0fffdffff9fffffffffffffffffffffc0000000000000000000000ff00000fffc040fffffffffffffffffffffffe0000000000000000000000ff00000fffc00067fffffffffffffffffffffe0000000000000000000000ff00000ffee00007ffffffffffffffffffffff0000000000000000000000ff000007fe40000fffffffffffffffffffffff8000000000000000000000ff000007fe00003fffffffffffffffffffffff8000000000000000000000ff00000fff00007fffffffffffffffffffffffc000000000000000000000ff000007ff0000fffffffffffffffffffffffff000000000000000000000ff00000fff0001fffffffffffffffffffffffff800000000000000000000;
assign cxk[2][32399:0] = 32400'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ff000000000000000000000000000000000000000000000000000000000fffe00000000000000000000000000000000000000000000000000000003fffff000000000000000000000000000000000000000000000000000000fffffff00000000000000000000000000000000000000000000000000001fffffffc0000000000000000000000000000000000000000000000000003fffffffe0000000000000000000000000000000000000000000000000007ffffffff000000000000000000000000000000000000000000000000000fffffffffc00000000000000000000000000000000000000000000000001fffffffffc00000000000000000000000000000000000000000000000003fffffffffe00000000000000000000000000000000000000000000000003ffffffffff00000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc000000000000000000000000000000000000000000000001fffffffffffc000000000000000000000000000000000000000000000007fffffffffffc00000000000000000000000000000000000000000000003ffffffffffff8000000000000000000000000000000000000000000007ffffffffffffff000000000000000000000000000000000000000000003ffffffffffffffe00000000000000000000000000000000000000000001fffffffffffffffc00000000000000000000000000000000000000000007fffffffffffffff80000000000000000000000000000000000000000001ffffffffffffffff0000000000000000000000000000000000000000001fffffffffffffffff000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000003ffffffffffffffffffc00000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffff80000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007fffffffffffffffffff8000000000000000000000000000000000000001ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000007ffffffffffffffffffffe000000000000000000000000000000000000007fffffffffffffffffffff00000000000000000000000000000000000001ffffffffffffffffffffff80000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000007ffffffffffffffffffffffe000000000000000000000000000000000000fffffffffffffffffffffffe000000000000000000000000000000000001ffffffffffffffffffffffff000000000000000000000000000000000007ffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffe0000000000000000000000000000000007ffffffffffffffffffffffffff000000000000000000000000000000000fffffffffffffffffffffffffff000000000000000000000000000000001fffffffffffffffffffffffffff800000000000000000000000000000003fffffffffffffffffffffffffff80000000000000000000000000000000ffffffffffffffffffffffffffffc0000000000000000000000000000001fffffe0fffffffffffffffffffff80000000000000000000000000000003fffffc07ffffffffffffffffffff80000000000000000000000000000007fffff807ffffffffffffffffffff8000000000000000000000000000000ffffff007ffffffffffffffffffff8000000000000000000000000000003ffffff003ffffffffffffffffffff8000000000000000000000000000007fffffe003ffffffffffffffffffff800000000000000000000000000000ffffffc003ffffffffffffffffffff800000000000000000000000000000ffffff0003ffffffffffffffffffff800000000000000000000000000001fffffe0003ffffffffffffffffffff800000000000000000000000000001fffffe0003ffffffffffffffffffff800000000000000000000000000003fffffe0003ffffffffffffffffffff800000000000000000000000000001fffffc0003ffffffffffffffffffff800000000000000000000000000001fffffc0007ffffffffffffffffffffc00000000000000000000000000000fffffc0007ffffffffffffffffffffc000000000000000000000000000003ffffc000fffffffffffffffffffffc000000000000000000000000000003ffffc000fffffffffffffffffffffe000000000000000000000000000001ffffc001fffffffffffffffffffffe000000000000000000000000000000ffffe003fffffffffffffffffffffe0000000000000000000000000000003ffff003ffffffffffffffffffffff0000000000000000000000000000000ffff80fffffffffffffffffffffff00000000000000000000000000000007ffffffffffffffffffffffffffff00000000000000000000000000000003ffffffffffffffffffffffffffff00000000000000000000000000000001ffffffffffffffffffffffffffff00000000000000000000000000000000ffffffffffffffffffffffffffff000000000000000000000000000000007fffffffffffffffffffffffffff000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000000ffffffffffffffffffffffffffe0000000000000000000000000000000007fffffffffffffffffffffffffe0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc00000000000000000000000000000000007ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff0000000000000000000000000000000000003fffffffffffffffffffffff0000000000000000000000000000000000001ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffff8000000000000000000ff000000e0000001ff83fffffffffffffffffffff8000000000000000000ff000001ff000001ff83fffffffffffffffffffff0000000000000000000ff000003fff80001ff87fffffffffffffffffffff0000000000000000000ff000007fff80001ff9fffffffffffffffffffffe0000000000000000000ff000007fffc0001ffffffffffffffffffffffffc0000000000000000000ff00000ffff00001ffffffffffffffffffffffff80000000000000000000ff00001ffff00001fffffffffffffffffffffffe00000000000000000000ff00000fffe00001fffffffffffffffffffffe0000000000000000000000ff000007ffc00001fffffffffffffffffffff80000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000003ff800001fffffffffffffffffffff00000000000000000000000ff000000fe000001fffffffffffffffffffff00000000000000000000000ff0e0000fc000001fffffffffffffffffffff00000000000000000000000ff3f800fff800601fffffffffffffffffffff80000000000000000000000ffffc00fffc03f01fffffffffffffffffffff80000000000000000000000fffff01fffe0ff81fffffffffffffffffffff80000000000000000000000ffffffffffffffc1fffffffffffffffffffffc0000000000000000000000ffcbffdfffffffe1fffffffffffffffffffffc0000000000000000000000ff819f0ffffffff9fffffffffffffffffffffc0000000000000000000000ff00040fffcc60fffffffffffffffffffffffe0000000000000000000000ff00000fffc0007ffffffffffffffffffffffe0000000000000000000000ff00000fffe0000fffffffffffffffffffffff0000000000000000000000ff000007fec0003fffffffffffffffffffffff0000000000000000000000ff000003fe00007fffffffffffffffffffffff8000000000000000000000ff000007ff0000ffffffffffffffffffffffffe000000000000000000000ff000007ff0001fffffffffffffffffffffffff000000000000000000000ff000007ff0003fffffffffffffffffffffffff800000000000000000000;
assign cxk[3][32399:0] = 32400'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ff000000000000000000000000000000000000000000000000000000000fffc00000000000000000000000000000000000000000000000000000003fffff000000000000000000000000000000000000000000000000000000fffffff00000000000000000000000000000000000000000000000000001fffffffc0000000000000000000000000000000000000000000000000003fffffffe0000000000000000000000000000000000000000000000000007ffffffff000000000000000000000000000000000000000000000000000fffffffffc00000000000000000000000000000000000000000000000001fffffffffc00000000000000000000000000000000000000000000000003fffffffffe00000000000000000000000000000000000000000000000003ffffffffff00000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc000000000000000000000000000000000000000000000000fffffffffffc000000000000000000000000000000000000000000000001fffffffffffc000000000000000000000000000000000000000000000007fffffffffffc00000000000000000000000000000000000000000000003ffffffffffff8000000000000000000000000000000000000000000007ffffffffffffff000000000000000000000000000000000000000000003ffffffffffffffe00000000000000000000000000000000000000000001fffffffffffffffc00000000000000000000000000000000000000000007fffffffffffffff80000000000000000000000000000000000000000001ffffffffffffffff0000000000000000000000000000000000000000001fffffffffffffffff000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000003ffffffffffffffffffc00000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffff80000000000000000000000000000000000000003fffffffffffffffffff8000000000000000000000000000000000000000ffffffffffffffffffff8000000000000000000000000000000000000001ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000007ffffffffffffffffffffe00000000000000000000000000000000000000ffffffffffffffffffffff00000000000000000000000000000000000001ffffffffffffffffffffff80000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000007ffffffffffffffffffffffe000000000000000000000000000000000000fffffffffffffffffffffffe000000000000000000000000000000000001ffffffffffffffffffffffff000000000000000000000000000000000007ffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffe0000000000000000000000000000000007ffffffffffffffffffffffffff000000000000000000000000000000000fffffffffffffffffffffffffff000000000000000000000000000000001fffffffffffffffffffffffffff800000000000000000000000000000003fffffffffffffffffffffffffff80000000000000000000000000000000ffffffffffffffffffffffffffffc0000000000000000000000000000001fffffe0fffffffffffffffffffff80000000000000000000000000000003fffffc07ffffffffffffffffffff80000000000000000000000000000007fffff807ffffffffffffffffffff8000000000000000000000000000000ffffff007ffffffffffffffffffff8000000000000000000000000000003ffffff003ffffffffffffffffffff8000000000000000000000000000007fffffe003ffffffffffffffffffff800000000000000000000000000000ffffffc003ffffffffffffffffffff800000000000000000000000000000ffffff0003ffffffffffffffffffff800000000000000000000000000001fffffe0003ffffffffffffffffffff800000000000000000000000000001fffffe0003ffffffffffffffffffff800000000000000000000000000003fffffe0003ffffffffffffffffffff800000000000000000000000000001fffffc0003ffffffffffffffffffff800000000000000000000000000001fffffc0007ffffffffffffffffffffc00000000000000000000000000000fffffc0007ffffffffffffffffffffc000000000000000000000000000003ffffc000fffffffffffffffffffffc000000000000000000000000000003ffffc000fffffffffffffffffffffe000000000000000000000000000001ffffc001fffffffffffffffffffffe000000000000000000000000000000ffffe003fffffffffffffffffffffe0000000000000000000000000000003ffff003ffffffffffffffffffffff0000000000000000000000000000000ffff80fffffffffffffffffffffff00000000000000000000000000000007ffffffffffffffffffffffffffff00000000000000000000000000000003ffffffffffffffffffffffffffff00000000000000000000000000000001ffffffffffffffffffffffffffff00000000000000000000000000000000ffffffffffffffffffffffffffff000000000000000000000000000000007fffffffffffffffffffffffffff000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000000ffffffffffffffffffffffffffe0000000000000000000000000000000007fffffffffffffffffffffffffe0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc00000000000000000000000000000000007ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff0000000000000000000000000000000000003fffffffffffffffffffffff0000000000000000000000000000000000000ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffff8000000000000000000ff000000f0000001ff83fffffffffffffffffffff8000000000000000000ff000001ff000001ff83fffffffffffffffffffff0000000000000000000ff000003fff80001ff87fffffffffffffffffffff0000000000000000000ff000007fff80001ff9fffffffffffffffffffffe0000000000000000000ff000007fffc0001ffffffffffffffffffffffffc0000000000000000000ff00000ffff00001ffffffffffffffffffffffff80000000000000000000ff00001ffff00001fffffffffffffffffffffffe00000000000000000000ff00000fffe00001fffffffffffffffffffffe0000000000000000000000ff000007ffc00001fffffffffffffffffffff80000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000003ff800001fffffffffffffffffffff00000000000000000000000ff000000fe000001fffffffffffffffffffff00000000000000000000000ff0e0000fc000001fffffffffffffffffffff00000000000000000000000ff3f800fff800601fffffffffffffffffffff80000000000000000000000ffffc00fffc03f01fffffffffffffffffffff80000000000000000000000fffff01fffe0ff81fffffffffffffffffffff80000000000000000000000ffffffffffffffc1fffffffffffffffffffffc0000000000000000000000ffcbffdfffffffe1fffffffffffffffffffffc0000000000000000000000ff819f0ffffffff9fffffffffffffffffffffc0000000000000000000000ff00040fffcc60fffffffffffffffffffffffe0000000000000000000000ff00000fffc0007ffffffffffffffffffffffe0000000000000000000000ff00000fffe0000fffffffffffffffffffffff0000000000000000000000ff000007fec0003fffffffffffffffffffffff0000000000000000000000ff000003fe00007fffffffffffffffffffffff8000000000000000000000ff000007ff0000ffffffffffffffffffffffffe000000000000000000000ff000007ff0001fffffffffffffffffffffffff000000000000000000000ff000007ff0003fffffffffffffffffffffffff800000000000000000000;
assign cxk[4][32399:0] = 32400'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fe000000000000000000000000000000000000000000000000000000000fffc00000000000000000000000000000000000000000000000000000003ffffe000000000000000000000000000000000000000000000000000000fffffff00000000000000000000000000000000000000000000000000001fffffff80000000000000000000000000000000000000000000000000003fffffffe0000000000000000000000000000000000000000000000000007ffffffff000000000000000000000000000000000000000000000000000fffffffff800000000000000000000000000000000000000000000000001fffffffffc00000000000000000000000000000000000000000000000003fffffffffe00000000000000000000000000000000000000000000000007ffffffffff00000000000000000000000000000000000000000000000007ffffffffff00000000000000000000000000000000000000000000000007ffffffffff00000000000000000000000000000000000000000000000007ffffffffff80000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffc000000000000000000000000000000000000000000000000fffffffffffc000000000000000000000000000000000000000000000001fffffffffff8000000000000000000000000000000000000000000000007fffffffffff800000000000000000000000000000000000000000000003ffffffffffff8000000000000000000000000000000000000000000007ffffffffffffff000000000000000000000000000000000000000000003ffffffffffffffe00000000000000000000000000000000000000000001fffffffffffffffc00000000000000000000000000000000000000000007fffffffffffffff00000000000000000000000000000000000000000001ffffffffffffffff0000000000000000000000000000000000000000001ffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000003ffffffffffffffffffc00000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000001fffffffffffffffffff80000000000000000000000000000000000000003fffffffffffffffffff8000000000000000000000000000000000000000ffffffffffffffffffff8000000000000000000000000000000000000001ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000007ffffffffffffffffffffe00000000000000000000000000000000000000ffffffffffffffffffffff00000000000000000000000000000000000001ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff80000000000000000000000000000000000007ffffffffffffffffffffffc000000000000000000000000000000000000fffffffffffffffffffffffe000000000000000000000000000000000003ffffffffffffffffffffffff000000000000000000000000000000000007ffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffe0000000000000000000000000000000007fffffffffffffffffffffffffe000000000000000000000000000000000fffffffffffffffffffffffffff000000000000000000000000000000001fffffffffffffffffffffffffff000000000000000000000000000000007fffffffffffffffffffffffffff80000000000000000000000000000000ffffffffffffffffffffffffffff80000000000000000000000000000001fffffe0fffffffffffffffffffff80000000000000000000000000000003fffffc07ffffffffffffffffffff00000000000000000000000000000007fffff807ffffffffffffffffffff0000000000000000000000000000001ffffff007ffffffffffffffffffff0000000000000000000000000000003ffffff003ffffffffffffffffffff0000000000000000000000000000007fffffc003ffffffffffffffffffff000000000000000000000000000000ffffff8003ffffffffffffffffffff000000000000000000000000000001ffffff0003ffffffffffffffffffff000000000000000000000000000001fffffe0003ffffffffffffffffffff000000000000000000000000000001fffffe0003ffffffffffffffffffff000000000000000000000000000001fffffe0003ffffffffffffffffffff000000000000000000000000000001fffffc0007ffffffffffffffffffff800000000000000000000000000001fffffc0007ffffffffffffffffffff8000000000000000000000000000007ffffc000fffffffffffffffffffffc000000000000000000000000000003ffffc000fffffffffffffffffffffc000000000000000000000000000003ffffc001fffffffffffffffffffffe000000000000000000000000000000ffffe001fffffffffffffffffffffe0000000000000000000000000000007fffe003fffffffffffffffffffffe0000000000000000000000000000003ffff007fffffffffffffffffffffe0000000000000000000000000000000ffffc0ffffffffffffffffffffffe00000000000000000000000000000007fffffffffffffffffffffffffffe00000000000000000000000000000003fffffffffffffffffffffffffffe00000000000000000000000000000001fffffffffffffffffffffffffffe000000000000000000000000000000007ffffffffffffffffffffffffffe000000000000000000000000000000003ffffffffffffffffffffffffffe000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000000ffffffffffffffffffffffffffe0000000000000000000000000000000007fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff0000000000000000000000000000000000007ffffffffffffffffffffffe0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000000ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffc00000000000000000000000000000000000007fffffffffffffffffffffc000000000000000000ff00000000000001ff83fffffffffffffffffffff8000000000000000000ff00000000000001ff83fffffffffffffffffffff8000000000000000000ff00000000000001ff83fffffffffffffffffffff8000000000000000000ff00000000000001ff83fffffffffffffffffffff0000000000000000000ff000000f0000001ff83fffffffffffffffffffff0000000000000000000ff000001ff000001ff87fffffffffffffffffffff0000000000000000000ff000003fff80001ff8fffffffffffffffffffffe0000000000000000000ff000007fff80001ffbfffffffffffffffffffffc0000000000000000000ff000007fffc0001ffffffffffffffffffffffff80000000000000000000ff00000ffff00001ffffffffffffffffffffffff00000000000000000000ff00001ffff00001fffffffffffffffffffffff800000000000000000000ff00000fffe00001fffffffffffffffffffffc0000000000000000000000ff000007ffc00001fffffffffffffffffffff00000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000003ff800001fffffffffffffffffffff00000000000000000000000ff000000fe000001fffffffffffffffffffff00000000000000000000000ff0e0000fc000001fffffffffffffffffffff00000000000000000000000ff3f800fff800601fffffffffffffffffffff00000000000000000000000ffffc00fffc03f01fffffffffffffffffffff80000000000000000000000fffff01fffe0ff81fffffffffffffffffffff80000000000000000000000ffffffffffffffc1fffffffffffffffffffff80000000000000000000000ffcbffdfffffffe1fffffffffffffffffffff80000000000000000000000ff819f0ffffffff1fffffffffffffffffffffc0000000000000000000000ff00040fffcc60fffffffffffffffffffffffc0000000000000000000000ff00000fffc0007ffffffffffffffffffffffe0000000000000000000000ff00000fffe0001ffffffffffffffffffffffe0000000000000000000000ff000007fec0003fffffffffffffffffffffff0000000000000000000000ff000003fe00007fffffffffffffffffffffffc000000000000000000000ff000007ff0000ffffffffffffffffffffffffe000000000000000000000ff000007ff0003fffffffffffffffffffffffff000000000000000000000ff000007ff0007fffffffffffffffffffffffff800000000000000000000;
assign cxk[5][32399:0] = 32400'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fff00000000000000000000000000000000000000000000000000000003fffffe00000000000000000000000000000000000000000000000000000fffffff80000000000000000000000000000000000000000000000000003fffffffe0000000000000000000000000000000000000000000000000007ffffffff800000000000000000000000000000000000000000000000000fffffffffc00000000000000000000000000000000000000000000000001ffffffffff00000000000000000000000000000000000000000000000003ffffffffff80000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffe000000000000000000000000000000000000000000000000ffffffffffff000000000000000000000000000000000000000000000000ffffffffffff000000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff8000000000000000000000000000000000000000003fff01ffffffffffff000000000000000000000000000000000000000001fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffc00000000000000000000000000000000000000001fffffffffffffffff8000000000000000000000000000000000000000003fffffffffffffffff000000000000000000000000000000000000000000ffffffffffffffffff000000000000000000000000000000000000000003fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff000000000000000000000000000000000000000007ffffffffffffffffff00000000000000000000000000000000000000000ffffffffffffffffffe00000000000000000000000000000000000000001ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffff80000000000000000000000000000000000000001fffffffffffffffffff80000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007fffffffffffffffffff8000000000000000000000000000000000000000ffffffffffffffffffffc000000000000000000000000000000000000001ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffe000000000000000000000000000000000000007ffffffffffffffffffffe00000000000000000000000000000000000000ffffffffffffffffffffff00000000000000000000000000000000000000ffffffffffffffffffffff80000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000003fffffffffffffffffffffff0000000000000000000000000000000000007fffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffffc00000000000000000000000000000000000ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffffe00000000000000000000000000000000003ffffffffffffffffffffffffe00000000000000000000000000000000007fffffffffffffffffffffffff00000000000000000000000000000000007ffffe0fffffffffffffffffff0000000000000000000000000000000000fffffe0fffffffffffffffffff0000000000000000000000000000000001fffffc0fffffffffffffffffff0000000000000000000000000000000001fffffc0fffffffffffffffffff8000000000000000000000000000000003fffffc0fffffffffffffffffff8000000000000000000000000000000003fffffc0fffffffffffffffffff8000000000000000000000000000000007fffffe1fffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff800000000000000000000000000000000fffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffffc000000000000000000000000000000003ffffffffffffffffffffffffffc000000000000000000000000000000003ffffffffffffffffffffffffffc000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000000fffffffffffffffffffffffffff0000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000003ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffffc00000000000000000000000000000000000ffffffffffffffffffffffffc000000000000000000000000000000000007fffffffffffffffffffffffe000000000000000000000000000000000007fffffffffffffffffffffffe000000000000000000000000000000000001fffffffffffffffffffffffe000000000000000000000000000000000000fffffffffffffffffffffffe0000000000000000000000000000000000007ffffffffffffffffffffffc0000000000000000000000000000000000003ffffffffffffffffffffffc0000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000000ffffffffffffffffffffff800000000000000000000000000000000000003fffffffffffffffffffff800000000000000000000000000000000000001fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff000000000000000000000000000000000000000fffffffffffffffffffff00000000000000000000ff00000000000001ff9fffffffffffffffffffff00000000000000000000ff00000000000001fffffffffffffffffffffffe00000000000000000000ff00000000000001fffffffffffffffffffffffc00000000000000000000ff00000000000001fffffffffffffffffffffffc00000000000000000000ff000000fe000001fffffffffffffffffffffff000000000000000000000ff000001ff800001ffffffffffffffffffffffc000000000000000000000ff000003fff80001fffffffffffffffffffff00000000000000000000000ff000003fff80001ffffffffffffffffffffe00000000000000000000000ff000003fffc0001ffffffffffffffffffffe00000000000000000000000ff000007fff00001ffffffffffffffffffffe00000000000000000000000ff00000ffff00001ffffffffffffffffffffe00000000000000000000000ff000007ffe00001ffffffffffffffffffffe00000000000000000000000ff000007ffc00001fffffffffffffffffffff00000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000001ff800001fffffffffffffffffffff00000000000000000000000ff0400007e000001fffffffffffffffffffff00000000000000000000000ff0f0001fe000001fffffffffffffffffffff00000000000000000000000ff1fc00fffc00701fffffffffffffffffffff00000000000000000000000ffffe00fffe03f81fffffffffffffffffffff80000000000000000000000fffffc1ffff0ffc1fffffffffffffffffffffc0000000000000000000000ffffffffffffffe1fffffffffffffffffffffe0000000000000000000000ffe1ffcffffffff3fffffffffffffffffffffe0000000000000000000000ffc08f0fffefffffffffffffffffffffffffff0000000000000000000000ff000007ffc0207fffffffffffffffffffffffc000000000000000000000ff00000fffc0003fffffffffffffffffffffffe000000000000000000000ff00000fffe0003ffffffffffffffffffffffff000000000000000000000ff000007ffc0003ffffffffffffffffffffffff800000000000000000000ff000003ff00007ffffffffffffffffffffffffc00000000000000000000ff000007ff8000ffffffffffffffffffffffffff00000000000000000000ff000003ff8001ffffffffffffffffffffffffff00000000000000000000ff000007ff8001ffffffffffffffffffffffffff00000000000000000000;
assign cxk[6][32399:0] = 32400'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003fff00000000000000000000000000000000000000000000000000000003fffffe00000000000000000000000000000000000000000000000000000fffffff80000000000000000000000000000000000000000000000000003fffffffe0000000000000000000000000000000000000000000000000007ffffffff800000000000000000000000000000000000000000000000000fffffffffc00000000000000000000000000000000000000000000000001ffffffffff00000000000000000000000000000000000000000000000003ffffffffff80000000000000000000000000000000000000000000000007ffffffffffc0000000000000000000000000000000000000000000000007ffffffffffe000000000000000000000000000000000000000000000000ffffffffffff000000000000000000000000000000000000000000000000ffffffffffff000000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff800000000000000000000000000000000000000000000001ffffffffffff8000000000000000000000000000000000000000003fff01ffffffffffff000000000000000000000000000000000000000001fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffc00000000000000000000000000000000000000001fffffffffffffffff8000000000000000000000000000000000000000003fffffffffffffffff000000000000000000000000000000000000000000ffffffffffffffffff000000000000000000000000000000000000000003fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff000000000000000000000000000000000000000007ffffffffffffffffff00000000000000000000000000000000000000000ffffffffffffffffffe00000000000000000000000000000000000000001ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffff80000000000000000000000000000000000000001fffffffffffffffffff80000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007fffffffffffffffffff8000000000000000000000000000000000000000ffffffffffffffffffffc000000000000000000000000000000000000001ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffe000000000000000000000000000000000000007ffffffffffffffffffffe00000000000000000000000000000000000000ffffffffffffffffffffff00000000000000000000000000000000000000ffffffffffffffffffffff80000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000003fffffffffffffffffffffff0000000000000000000000000000000000007fffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffffc00000000000000000000000000000000000ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffffe00000000000000000000000000000000003ffffffffffffffffffffffffe00000000000000000000000000000000007fffffffffffffffffffffffff00000000000000000000000000000000007ffffe0fffffffffffffffffff0000000000000000000000000000000000fffffe0fffffffffffffffffff0000000000000000000000000000000001fffffc0fffffffffffffffffff0000000000000000000000000000000001fffffc0fffffffffffffffffff8000000000000000000000000000000003fffffc0fffffffffffffffffff8000000000000000000000000000000003fffffc0fffffffffffffffffff8000000000000000000000000000000007fffffe1fffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff800000000000000000000000000000000fffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000007ffffffffffffffffffffffffffc000000000000000000000000000000003ffffffffffffffffffffffffffc000000000000000000000000000000003ffffffffffffffffffffffffffc000000000000000000000000000000001ffffffffffffffffffffffffffe000000000000000000000000000000000fffffffffffffffffffffffffff0000000000000000000000000000000007ffffffffffffffffffffffffff8000000000000000000000000000000003ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc0000000000000000000000000000000000fffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000001ffffffffffffffffffffffffc00000000000000000000000000000000000ffffffffffffffffffffffffc000000000000000000000000000000000007fffffffffffffffffffffffe000000000000000000000000000000000007fffffffffffffffffffffffe000000000000000000000000000000000001fffffffffffffffffffffffe000000000000000000000000000000000000fffffffffffffffffffffffe0000000000000000000000000000000000007ffffffffffffffffffffffc0000000000000000000000000000000000003ffffffffffffffffffffffc0000000000000000000000000000000000001ffffffffffffffffffffffc0000000000000000000000000000000000000ffffffffffffffffffffff800000000000000000000000000000000000003fffffffffffffffffffff800000000000000000000000000000000000001fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffff000000000000000000000000000000000000000fffffffffffffffffffff00000000000000000000ff00000000000001ff9fffffffffffffffffffff00000000000000000000ff00000000000001fffffffffffffffffffffffe00000000000000000000ff00000000000001fffffffffffffffffffffffc00000000000000000000ff00000000000001fffffffffffffffffffffffc00000000000000000000ff000000fe000001fffffffffffffffffffffff000000000000000000000ff000001ff800001ffffffffffffffffffffffc000000000000000000000ff000003fff80001fffffffffffffffffffff00000000000000000000000ff000003fff80001ffffffffffffffffffffe00000000000000000000000ff000003fffc0001ffffffffffffffffffffe00000000000000000000000ff00000ffff00001ffffffffffffffffffffe00000000000000000000000ff00000ffff00001ffffffffffffffffffffe00000000000000000000000ff000007ffe00001ffffffffffffffffffffe00000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000007ff800001fffffffffffffffffffff00000000000000000000000ff000001ff800001fffffffffffffffffffff00000000000000000000000ff0400007e000001fffffffffffffffffffff00000000000000000000000ff0f0003fe000001fffffffffffffffffffff00000000000000000000000ff1fc00fffc00701fffffffffffffffffffff00000000000000000000000ffbfe00fffe03f81fffffffffffffffffffff80000000000000000000000fffff81ffff0ffc1fffffffffffffffffffffc0000000000000000000000ffffffffffffffe1fffffffffffffffffffffe0000000000000000000000ffe1ffcffffffff3fffffffffffffffffffffe0000000000000000000000ffc08f0fffefffffffffffffffffffffffffff0000000000000000000000ff000007ffc0207fffffffffffffffffffffffc000000000000000000000ff00000fffc0003fffffffffffffffffffffffe000000000000000000000ff00000fffe0001ffffffffffffffffffffffff000000000000000000000ff000007ffc0003ffffffffffffffffffffffff800000000000000000000ff000003ff00007ffffffffffffffffffffffffc00000000000000000000ff000007ff8000ffffffffffffffffffffffffff00000000000000000000ff000003ff8001ffffffffffffffffffffffffff00000000000000000000ff000007ff8001ffffffffffffffffffffffffff00000000000000000000;
assign cxk[7][32399:0] = 32400'h000000000000000000000000000001ffffffffffc0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003fffffffffff0000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000003800007fffffffffff800000000000000000000000000000000000000003fffc007fffffffffff00000000000000000000000000000000000000000fffff00fffffffffffe00000000000000000000000000000000000000003fffffffffffffffff000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000000000000000000003fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffff800000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffffc0000000000000000000000000000000000000001fffffffffffffffffffc0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000007ffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffffc00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000001ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff80000000000000000000000000000000000007ffffffffffffffffffffff8000000000000000000000000000000000000fffffffffffffffffffffffc000000000000000000000000000000000001fffffffffffffffffffffffe000000000000000000000000000000000001ffffffffffffffffffffffff000000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000007ffffffffffffffffffffffffe00000000000000000000000000000000007ffffffffffffffffffffffffe0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffe0000000000000000000000000000000000fffffffffffffffffffffffffe00000000000000000000000000000000007fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000001fffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffff800000000000000000000000000000000007ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff8000000000000000000000000000000000007fffffffffffffffffffffff0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000001ffffffffffffffffffffffe0000000000000000000000000000000000000ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000000fffffffffffffffffffffe000000000000000000000000000000000000007ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffff0000000000000000000000000000000000000000003ffffffffffffffffe000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff000000fe000001ffffffffffffffffffff000000000000000000000000ff000001ff800001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff800000000000000000000000ff000003fffc0001ffffffffffffffffffff800000000000000000000000ff00000ffff00001ffffffffffffffffffffc00000000000000000000000ff00000ffff00001ffffffffffffffffffffc00000000000000000000000ff000007ffe00001ffffffffffffffffffffc00000000000000000000000ff000007ff800001ffffffffffffffffffffe00000000000000000000000ff000007ff800001ffffffffffffffffffffe00000000000000000000000ff000001ff800001fffffffffffffffffffff00000000000000000000000ff0400007e000001fffffffffffffffffffff00000000000000000000000ff0f0003fe000001fffffffffffffffffffff00000000000000000000000ff1fc00fffc00701fffffffffffffffffffff80000000000000000000000ffbfe00fffe03f81fffffffffffffffffffffc0000000000000000000000fffff81ffff0ffc1fffffffffffffffffffffe0000000000000000000000ffffffffffffffe3ffffffffffffffffffffff0000000000000000000000ffe1ffcffffffff3ffffffffffffffffffffff8000000000000000000000ffc08f0fffefffffffffffffffffffffffffff8000000000000000000000ff000007ffc0207fffffffffffffffffffffffc000000000000000000000ff00000fffc0003ffffffffffffffffffffffff000000000000000000000ff00000fffe0001ffffffffffffffffffffffff000000000000000000000ff000007ffc0003ffffffffffffffffffffffff800000000000000000000ff000003ff00007ffffffffffffffffffffffffc00000000000000000000ff000007ff8000fffffffffffffffffffffffffe00000000000000000000ff000003ff8000ffffffffffffffffffffffffff00000000000000000000ff000007ff8001ffffffffffffffffffffffffff00000000000000000000;
assign cxk[8][32399:0] = 32400'h000000000000000000000000000001ffffffffffc0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003fffffffffff0000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000003800007fffffffffff800000000000000000000000000000000000000003fffc007fffffffffff00000000000000000000000000000000000000000fffff00fffffffffffe00000000000000000000000000000000000000003fffffffffffffffff000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000000000000000000003fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffff800000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffffc0000000000000000000000000000000000000001fffffffffffffffffffc0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000007ffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffffc00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000001ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff80000000000000000000000000000000000007ffffffffffffffffffffff8000000000000000000000000000000000000fffffffffffffffffffffffc000000000000000000000000000000000001fffffffffffffffffffffffe000000000000000000000000000000000001ffffffffffffffffffffffff000000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000007ffffffffffffffffffffffffe00000000000000000000000000000000007ffffffffffffffffffffffffe0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffe0000000000000000000000000000000000fffffffffffffffffffffffffe00000000000000000000000000000000007fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000001fffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffff800000000000000000000000000000000007ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff8000000000000000000000000000000000007fffffffffffffffffffffff0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000001ffffffffffffffffffffffe0000000000000000000000000000000000000ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000000fffffffffffffffffffffe000000000000000000000000000000000000007ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffff0000000000000000000000000000000000000000003ffffffffffffffffe000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff000000fe000001ffffffffffffffffffff000000000000000000000000ff000001ff800001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff800000000000000000000000ff000003fffc0001ffffffffffffffffffff800000000000000000000000ff000007fff00001ffffffffffffffffffffc00000000000000000000000ff00000ffff00001ffffffffffffffffffffc00000000000000000000000ff000007ffe00001ffffffffffffffffffffc00000000000000000000000ff000007ff800001ffffffffffffffffffffe00000000000000000000000ff000007ff800001ffffffffffffffffffffe00000000000000000000000ff000001ff800001fffffffffffffffffffff00000000000000000000000ff0400007c000001fffffffffffffffffffff00000000000000000000000ff0f0001fe000001fffffffffffffffffffff00000000000000000000000ff1fc00fffc00701fffffffffffffffffffff80000000000000000000000ffbfe00fffe03f81fffffffffffffffffffffc0000000000000000000000fffffc1ffff0ffc1fffffffffffffffffffffe0000000000000000000000ffffffffffffffe3ffffffffffffffffffffff0000000000000000000000ffe1ffcffffffff3ffffffffffffffffffffff8000000000000000000000ffc08f0fffefffffffffffffffffffffffffff8000000000000000000000ff000007ffc0207fffffffffffffffffffffffc000000000000000000000ff00000fffc0003ffffffffffffffffffffffff000000000000000000000ff00000fffe0001ffffffffffffffffffffffff000000000000000000000ff000007ffc0003ffffffffffffffffffffffff800000000000000000000ff000003ff00007ffffffffffffffffffffffffc00000000000000000000ff000007ff8000fffffffffffffffffffffffffe00000000000000000000ff000003ff8000ffffffffffffffffffffffffff00000000000000000000ff000007ff8001ffffffffffffffffffffffffff00000000000000000000;
assign cxk[9][32399:0] = 32400'h000000000000000000000000000001ffffffffffc0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003ffffffffffe0000000000000000000000000000000000000000000000003fffffffffff0000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff0000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000000000007fffffffffff8000000000000000000000000000000000000000003800007fffffffffff800000000000000000000000000000000000000003fffc007fffffffffff00000000000000000000000000000000000000000fffff00fffffffffffe00000000000000000000000000000000000000003fffffffffffffffff000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000000000000000000003fffffffffffffffffe000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff000000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000001ffffffffffffffffffc00000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007fffffffffffffffffe00000000000000000000000000000000000000000ffffffffffffffffffc00000000000000000000000000000000000000000ffffffffffffffffff800000000000000000000000000000000000000001ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000003ffffffffffffffffff800000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffffffc0000000000000000000000000000000000000001fffffffffffffffffffc0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000007ffffffffffffffffffff800000000000000000000000000000000000000fffffffffffffffffffffc00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000001ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff00000000000000000000000000000000000003ffffffffffffffffffffff80000000000000000000000000000000000007ffffffffffffffffffffff8000000000000000000000000000000000000fffffffffffffffffffffffc000000000000000000000000000000000001fffffffffffffffffffffffe000000000000000000000000000000000001ffffffffffffffffffffffff000000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000003ffffffffffffffffffffffffc00000000000000000000000000000000007ffffffffffffffffffffffffe00000000000000000000000000000000007ffffffffffffffffffffffffe0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000000ffffffffffffffffffffffffff0000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000001ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff8000000000000000000000000000000000ffffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffff80000000000000000000000000000000007fffffffffffffffffffffffffc0000000000000000000000000000000003fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffc0000000000000000000000000000000001fffffffffffffffffffffffffe0000000000000000000000000000000000fffffffffffffffffffffffffe00000000000000000000000000000000007fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000003fffffffffffffffffffffffff00000000000000000000000000000000001fffffffffffffffffffffffff80000000000000000000000000000000000fffffffffffffffffffffffff800000000000000000000000000000000007ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000003ffffffffffffffffffffffff800000000000000000000000000000000001ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff800000000000000000000000000000000000ffffffffffffffffffffffff8000000000000000000000000000000000007fffffffffffffffffffffff0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000003ffffffffffffffffffffffe0000000000000000000000000000000000001ffffffffffffffffffffffe0000000000000000000000000000000000000ffffffffffffffffffffffe00000000000000000000000000000000000007fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000003fffffffffffffffffffffe00000000000000000000000000000000000001fffffffffffffffffffffe00000000000000000000000000000000000000fffffffffffffffffffffe000000000000000000000000000000000000007ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffffc000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff8000000000000000000000000000000000000003ffffffffffffffffffff0000000000000000000000000000000000000003fffffffffffffffffffe0000000000000000000000000000000000000003fffffffffffffffffff80000000000000000000000000000000000000007ffffffffffffffffff80000000000000000000000000000000000000000fffffffffffffffff0000000000000000000000000000000000000000003ffffffffffffffffe000000000000000000000000000000000000000000fffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff00000000000001fffffffffffffffffffe000000000000000000000000ff000001ff000001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff000000000000000000000000ff000003fff80001ffffffffffffffffffff000000000000000000000000ff000003fffc0001ffffffffffffffffffff800000000000000000000000ff000003fff80001ffffffffffffffffffff800000000000000000000000ff00000ffff00001ffffffffffffffffffffc00000000000000000000000ff00000fffe00001ffffffffffffffffffffc00000000000000000000000ff000003ffc00001ffffffffffffffffffffc00000000000000000000000ff000003ffc00001ffffffffffffffffffffe00000000000000000000000ff000003ffc00001ffffffffffffffffffffe00000000000000000000000ff000000ff000001fffffffffffffffffffff00000000000000000000000ff0300007e000001fffffffffffffffffffff00000000000000000000000ff07c007ffc00181fffffffffffffffffffff00000000000000000000000ff0ff007ffe00fc1fffffffffffffffffffff80000000000000000000000ff3ffc0ffff03fc1fffffffffffffffffffffc0000000000000000000000ffffffffffffffe1fffffffffffffffffffffe0000000000000000000000fffffffffffffffbffffffffffffffffffffff0000000000000000000000fff07fcfffffffffffffffffffffffffffffff8000000000000000000000ff000307ffe3183fffffffffffffffffffffff8000000000000000000000ff000007ffe0003fffffffffffffffffffffffc000000000000000000000ff000007ffe0001ffffffffffffffffffffffff000000000000000000000ff000007ffe0001ffffffffffffffffffffffff000000000000000000000ff000001ff80003ffffffffffffffffffffffff800000000000000000000ff000001ff80007ffffffffffffffffffffffffc00000000000000000000ff000003ffc000fffffffffffffffffffffffffe00000000000000000000ff000003ffc000ffffffffffffffffffffffffff00000000000000000000ff000003ffc001ffffffffffffffffffffffffff00000000000000000000;
//assign cxk[0][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[1][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[2][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[3][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[4][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[5][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[6][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[7][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[8][32399:0] = 32400'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//assign cxk[9][32399:0] = 32400'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000000000000000000000e00000000000000000000000000000000000000000000000000000000000e00000000000000000000000000000000000000000000000100000000000e00000000000000000000000000000000000000000000000100000004000f0000000000000000000000000000000000000000000000038000000c001f000000000000000000000000000000000000000000000007c000001f003f80000000000000000000000000000000000000000000001fffffffff807fc00000000000000000000000000000000000000000000007c018001e001f000000000000000000000000000000000000000000000007c03c000c000e000000000000000000000000000000000000000000000007c8182005cc041c0000000000000000000000000000000000000000000007dffff9ffcfffff0000000000000000000000000000000000000000000007df00fc1fef8e3f0000000000000000000000000000000000000000000007df0078cfef8e3e0000000000000000000000000000000000000000000007df0079ce0f9f3e0000000000000000000000000000000000000000000007dffe79ce0ffffe0000000000000000000000000000000000000000000007df0079ceeffffe0000000000000000000000000000000000000000000007df0079ceefbfbe0000000000000000000000000000000000000000000007df00f9ceef8e3e00000000000000000000000000000000000000000000079ffff9ceef8e3e00000000000000000000000000000000000000000000079c3c71ceeffffe0000000000000000000000000000000000000000000007803c01cecf863e0000000000000000000000000000000000000000000007073c71cecf041e000000000000000000000000000000000000000000000f3f3cfdde0e0e06000000000000000000000000000000000000000000000effbdffde001f00000000000000000000000000000000000000000000001cf83c0f9e007fe00000000000000000000000000000000000000000000038603c071e003f800000000000000000000000000000000000000000000020303c0c1e001f0000000000000000000000000000000000000000000000000038001c001f0000000000000000000000000000000000000000000000000038001c000e00000000000000000000000000000000000000000000000000200000000e00000000000000000000000000000000000000000000000000000000000e00000000000000000000000000000000000000000000000000000000000e000000000000000000000000000000000000000000000000000000000006000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040000000000000000000000000000000000000080000004000000000000040000000000000000000400000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000004008000400000000000000000000800000000000000000000000000000004008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000100000001000000000000000000000000000000000000000000000000000110000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
always@(posedge clk or negedge resetn) begin
	if (~resetn) begin
		clk_cnt <= 0;
		cmd_index <= 0;
		init_state <= INIT_RESET;
        
        time_cnt<= 4'b0000;
		lcd_cs_r <= 1;
		lcd_rs_r <= 1;
		lcd_reset_r <= 0;
		spi_data <= 8'hFF;
		bit_loop <= 0;

		pixel_cnt <= 0;
	end else begin

		case (init_state)

			INIT_RESET : begin
				if (clk_cnt == CNT_100MS) begin
					clk_cnt <= 0;
					init_state <= INIT_PREPARE;
					lcd_reset_r <= 1;
				end else begin
					clk_cnt <= clk_cnt + 1;
				end
			end

			INIT_PREPARE : begin
				if (clk_cnt == CNT_200MS) begin
					clk_cnt <= 0;
					init_state <= INIT_WAKEUP;
				end else begin
					clk_cnt <= clk_cnt + 1;
				end
			end

			INIT_WAKEUP : begin
				if (bit_loop == 0) begin
					// start
					lcd_cs_r <= 0;
					lcd_rs_r <= 0;
					spi_data <= 8'h11; // exit sleep
					bit_loop <= bit_loop + 1;
				end else if (bit_loop == 8) begin
					// end
					lcd_cs_r <= 1;
					lcd_rs_r <= 1;
					bit_loop <= 0;
					init_state <= INIT_SNOOZE;
				end else begin
					// loop
					spi_data <= { spi_data[6:0], 1'b1 };
					bit_loop <= bit_loop + 1;
				end
			end

			INIT_SNOOZE : begin
				if (clk_cnt == CNT_120MS) begin
					clk_cnt <= 0;
					init_state <= INIT_WORKING;
				end else begin
					clk_cnt <= clk_cnt + 1;
				end
			end

			INIT_WORKING : begin
				if (cmd_index == MAX_CMDS + 1) begin
					init_state <= INIT_DONE;
				end else begin
					if (bit_loop == 0) begin
						// start
						lcd_cs_r <= 0;
						lcd_rs_r <= init_cmd[cmd_index][8];
						spi_data <= init_cmd[cmd_index][7:0];
						bit_loop <= bit_loop + 1;
					end else if (bit_loop == 8) begin
						// end
						lcd_cs_r <= 1;
						lcd_rs_r <= 1;
						bit_loop <= 0;
						cmd_index <= cmd_index + 1; // next command
					end else begin
						// loop
						spi_data <= { spi_data[6:0], 1'b1 };
						bit_loop <= bit_loop + 1;
					end
				end
			end

			INIT_DONE : begin
                if(time_cnt == 10) begin
                    time_cnt<=4'b0000;
                end
				if (pixel_cnt == 32400) begin
					time_cnt<=time_cnt+1'b1;
                    pixel_cnt<=0;
				end else begin //一个像素点需要分上下两次来运，一次只能运8bit
					if (bit_loop == 0) begin
						// start
						lcd_cs_r <= 0;
						lcd_rs_r <= 1;
//						spi_data <= 8'hF8; // RED
                            if(cxk[time_cnt][pixel_cnt]==1'b1) begin 
                                spi_data <= 8'h00;
                            end
                            else begin
                                spi_data <= 8'hff;
                            end
						bit_loop <= bit_loop + 1;
					end else if (bit_loop == 8) begin
						// next byte
//						spi_data <= 8'h00; // RED
                            if(cxk[time_cnt][pixel_cnt]==1'b1) begin 
                                spi_data <= 8'h00;
                            end
                            else begin
                                spi_data <= 8'hff;
                            end
						bit_loop <= bit_loop + 1;
					end else if (bit_loop == 16) begin
						// end
						lcd_cs_r <= 1;
						lcd_rs_r <= 1;
						bit_loop <= 0;
						pixel_cnt <= pixel_cnt + 1; // next pixel
					end else begin
						// loop
						spi_data <= { spi_data[6:0], 1'b1 };
						bit_loop <= bit_loop + 1;
					end
				end
			end
		endcase

	end
end

endmodule
